-- EX Stage
-- Author:  Anshul Kharbanda
-- Created: 11 - 29 - 2018
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ex_stage is
    port (
        clk: in std_logic
    );
end entity;

architecture arch of ex_stage is
begin
    -- ALU
    -- Branch
    -- Forwarding
end architecture;
